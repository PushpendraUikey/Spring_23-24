*Zener Regulator
Vin Supply Gnd 0
*Series limiter
RS Supply Zplus 300
*Zener modeled as a diode with low breakdown voltage of 4.7V
D1 Ztest Zplus DF
.MODEL DF D (IS=6.22n N=1.9224 RS=0.336 CJ0=764f VJ=0.75 BV=4.7 TT=2.88n)
*0V source inserted to measure Zener current
VZtest Ztest Gnd 0
*Load resistor
RL Zplus Rtest 1000
*0V source inserted to measure current through the load resistor
VRtest Rtest Gnd 0
*DC analysis: Sweep input voltage
.DC Vin -2.0 12.0 0.05 
.control
run
plot V(Zplus) ylimit 0 5.5
plot I(VZtest) ylimit 0 5.5m
plot I(VRtest)
.endc
.end

